`include "define.v"

`resetall
`timescale 1ns / 1ps
`default_nettype none

module processor #(
  parameter [31:0] PC_BASE_ADDR = `CPU_PC_BASE_ADDR,
  parameter [31:0] SP_BASE_ADDR = `CPU_SP_BASE_ADDR
)(
  input         clk,
  input         rst,
  output [31:0] mem_addr_o,
  output        mem_rstrb_o,
  input  [31:0] mem_rdata_i,
  output [3:0]  mem_wmask_o,
  output [31:0] mem_wdata_o
);

// define register file
reg [31:0] regfile_ra[0:31];  // ra: reg array

// ----------------------------------------------------------------------------
// with reset the regfile is synthesized to SB_DFFESR and SB_LUT4
// ----------------------------------------------------------------------------
// genvar i;
// generate
//   for (i = 0; i < 31; i = i + 1) begin
//     always @(posedge clk) begin
//       if (rst) begin
//         regfile_ra[i] <= 32'b0;
//       end
//       else if ((wb_en_w) & (rd_id_w == (i))) begin
//         regfile_ra[i] <= wb_data_w;
//       end
//     end
//   end
// endgenerate

// ----------------------------------------------------------------------------
// with reset the regfile is synthesized to SB_DFFESR and SB_LUT4
// ----------------------------------------------------------------------------
// integer i;
// always @(posedge clk) begin
//   if (rst) begin
//     for (i = 0; i < 31; ++i) begin
//       regfile_ra[i] <= 32'b0;
//     end
//   end
//   else if (wb_en_w) begin
//     regfile_ra[rd_id_w] <= wb_data_w;
//   end
// end

// ----------------------------------------------------------------------------
// without reset the regfile is synthesized to SB_RAM40_4K
// ----------------------------------------------------------------------------
integer i;
initial begin
  for (i = 0; i < 32; i = i + 1) begin
    regfile_ra[i] = 0;
  end
  regfile_ra[`sp] = SP_BASE_ADDR;
end

always @(posedge clk) begin
  if (wb_en_w) begin
    regfile_ra[rd_id_w] <= wb_data_w;
  end
end

// ----------------------------------------------------------------------------
// CPU State Machine
// ----------------------------------------------------------------------------
// define state parameter
localparam IF  = 0;
localparam ID  = 1;
localparam EXE = 2;
localparam MEM = 3;
localparam WB  = 4;

reg [2:0] state_r;
always @(posedge clk) begin
  if (rst) begin
    state_r <= WB;
    inst_r <= 32'b0;
  end
  else begin
    case (state_r)
      IF: begin
        state_r <= ID;
        inst_r <= mem_rdata_i;
      end
      ID: begin
        state_r <= EXE;
      end
      EXE: begin
        if (is_load_w | is_store_w) begin
          state_r <= MEM;
        end
        else begin
          state_r <= WB;
        end
      end
      MEM: begin
        state_r <= WB;
      end
      WB: begin
        state_r <= IF;
      end
      default: begin
        state_r <= WB;
      end 
    endcase
  end
end

// ----------------------------------------------------------------------------
// Instruction Decoder
// ----------------------------------------------------------------------------
reg [31:0] inst_r;

wire is_alu_reg_w = inst_r[6:0] == 7'b011_0011;   // rd <- rs1 OP rs2
wire is_alu_imm_w = inst_r[6:0] == 7'b001_0011;   // rd <- rs1 OP Iimm
wire is_branch_w  = inst_r[6:0] == 7'b110_0011;   // if(rs1 OP rs2) PC <- PC + Bimm
wire is_jalr_w    = inst_r[6:0] == 7'b110_0111;   // rd <- PC + 4; PC <- rs1 + Iimm
wire is_jal_w     = inst_r[6:0] == 7'b110_1111;   // rd <- PC + 4; PC <- PC + Jimm
wire is_auipc_w   = inst_r[6:0] == 7'b001_0111;   // rd <- PC + Uimm
wire is_lui_w     = inst_r[6:0] == 7'b011_0111;   // rd <- Uimm
wire is_load_w    = inst_r[6:0] == 7'b000_0011;   // rd <- MEM[rs1 + Iimm]
wire is_store_w   = inst_r[6:0] == 7'b010_0011;   // MEM[rs1 + Simm] <- rs2
wire is_system_w  = inst_r[6:0] == 7'b111_0011;   // special

wire [4:0] rs1_id_w = inst_r[19:15];
wire [4:0] rs2_id_w = inst_r[24:20];
wire [4:0] rd_id_w  = inst_r[11:7];

reg [31:0] rs1_r;
reg [31:0] rs2_r;
always @(posedge clk) begin
  if (rst) begin
    rs1_r <= 32'b0;
    rs2_r <= 32'b0;
  end
  else if (state_r == ID) begin
    rs1_r <= regfile_ra[rs1_id_w];
    rs2_r <= regfile_ra[rs2_id_w];
  end
end

wire [2:0] funct3_w = inst_r[14:12];
wire [6:0] funct7_w = inst_r[31:25];

wire [31:0] Iimm_w = {{21{inst_r[31]}}, inst_r[30:20]};
wire [31:0] Uimm_w = {    inst_r[31],   inst_r[30:12], {12{1'b0}}};
wire [31:0] Simm_w = {{21{inst_r[31]}}, inst_r[30:25], inst_r[11:7]};
wire [31:0] Bimm_w = {{20{inst_r[31]}}, inst_r[7], inst_r[30:25], inst_r[11:8], 1'b0};
wire [31:0] Jimm_w = {{12{inst_r[31]}}, inst_r[19:12], inst_r[20], inst_r[30:21], 1'b0};

// ----------------------------------------------------------------------------
// Instruction Monitor (debug only)
// ----------------------------------------------------------------------------
always @(posedge clk) begin
  if (state_r == EXE) begin
    case (1'b1)
      is_alu_reg_w: begin
        // $display("[%t ps][CPU ]: rd[%d] <- rs1[%d] OP rs2[%d]", $realtime, rd_id_w, rs1_id_w, rs2_id_w);
        case (funct3_w)
          3'b000: begin
            if (funct7_w[5]) begin
              $display("[%t ps][CPU ]: SUB rd[%d], rs1[%d](%h), rs2[%d](%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, rs2_id_w, rs2_r);
            end
            else begin
              $display("[%t ps][CPU ]: ADD rd[%d], rs1[%d](%h), rs2[%d](%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, rs2_id_w, rs2_r);
            end
          end
          3'b001: $display("[%t ps][CPU ]: SLL rd[%d], rs1[%d](%h), rs2[%d](%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, rs2_id_w, rs2_r);
          3'b010: $display("[%t ps][CPU ]: SLT rd[%d], rs1[%d](%h), rs2[%d](%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, rs2_id_w, rs2_r);
          3'b011: $display("[%t ps][CPU ]: SLTU rd[%d], rs1[%d](%h), rs2[%d](%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, rs2_id_w, rs2_r);
          3'b100: $display("[%t ps][CPU ]: XOR rd[%d], rs1[%d](%h), rs2[%d](%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, rs2_id_w, rs2_r);
          3'b101: begin
            if (funct7_w[5]) begin
              $display("[%t ps][CPU ]: SRA rd[%d], rs1[%d](%h), rs2[%d](%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, rs2_id_w, rs2_r);
            end
            else begin
              $display("[%t ps][CPU ]: SRL rd[%d], rs1[%d](%h), rs2[%d](%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, rs2_id_w, rs2_r);
            end
          end
          3'b110: $display("[%t ps][CPU ]: OR rd[%d], rs1[%d](%h), rs2[%d](%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, rs2_id_w, rs2_r);
          3'b111: $display("[%t ps][CPU ]: AND rd[%d], rs1[%d](%h), rs2[%d](%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, rs2_id_w, rs2_r);
        endcase
      end
      is_alu_imm_w: begin
        // $display("[%t ps][CPU ]: rd[%d] <- rs1[%d] OP Iimm(%h)", $realtime, rd_id_w, rs1_id_w, Iimm_w);
        case (funct3_w)
          3'b000: $display("[%t ps][CPU ]: ADDI rd[%d], rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, Iimm_w);
          3'b001: $display("[%t ps][CPU ]: SLLI rd[%d], rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, Iimm_w);
          3'b010: $display("[%t ps][CPU ]: SLTI rd[%d], rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, Iimm_w);
          3'b011: $display("[%t ps][CPU ]: SLTUI rd[%d], rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, Iimm_w);
          3'b100: $display("[%t ps][CPU ]: XORI rd[%d], rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, Iimm_w);
          3'b101: begin
            if (funct7_w[5]) begin
              $display("[%t ps][CPU ]: SRAI rd[%d], rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, Iimm_w);
            end
            else begin
              $display("[%t ps][CPU ]: SRLI rd[%d], rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, Iimm_w);
            end
          end
          3'b110: $display("[%t ps][CPU ]: ORI rd[%d], rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, Iimm_w);
          3'b111: $display("[%t ps][CPU ]: ANDI rd[%d], rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, Iimm_w);
        endcase
      end
      is_branch_w: begin
        // $display("[%t ps][CPU ]: if(rs1[%d] OP rs2[%d]) PC <- PC(%d) + Bimm(%h)", $realtime, rs1_id_w, rs2_id_w, pc_r, Bimm_w);
        case (funct3_w)
          3'b000: $display("[%t ps][CPU ]: BEQ rs1[%d](%h), rs2[%d](%h), Bimm(%h)", $realtime, rs1_id_w, rs1_r, rs2_id_w, rs2_r, Bimm_w);
          3'b001: $display("[%t ps][CPU ]: BNE rs1[%d](%h), rs2[%d](%h), Bimm(%h)", $realtime, rs1_id_w, rs1_r, rs2_id_w, rs2_r, Bimm_w);
          3'b100: $display("[%t ps][CPU ]: BLT rs1[%d](%h), rs2[%d](%h), Bimm(%h)", $realtime, rs1_id_w, rs1_r, rs2_id_w, rs2_r, Bimm_w);
          3'b101: $display("[%t ps][CPU ]: BGE rs1[%d](%h), rs2[%d](%h), Bimm(%h)", $realtime, rs1_id_w, rs1_r, rs2_id_w, rs2_r, Bimm_w);
          3'b110: $display("[%t ps][CPU ]: BLTU rs1[%d](%h), rs2[%d](%h), Bimm(%h)", $realtime, rs1_id_w, rs1_r, rs2_id_w, rs2_r, Bimm_w);
          3'b111: $display("[%t ps][CPU ]: BGEU rs1[%d](%h), rs2[%d](%h), Bimm(%h)", $realtime, rs1_id_w, rs1_r, rs2_id_w, rs2_r, Bimm_w);
          default: $display("[%t ps][CPU ]: Wrong Branch, check funct3: x[%d](%h), x[%d](%h), Bimm(%h)", $realtime, rs1_id_w, rs1_r, rs2_id_w, rs2_r, Bimm_w);
        endcase
      end
      is_jalr_w: begin
        // $display("[%t ps][CPU ]: rd[%d] <- PC(%d) + 4; PC <- rs1[%d] + Iimm(%h)", $realtime, rd_id_w, pc_r, rs1_id_w, Iimm_w);
        $display("[%t ps][CPU ]: JALR rd[%d](%h), rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, (pc_r + 4), rs1_id_w, rs1_r, Iimm_w);
      end
      is_jal_w: begin
        // $display("[%t ps][CPU ]: rd[%d] <- PC(%d) + 4; PC <- PC + Jimm(%h)", $realtime, rd_id_w, pc_r, Jimm_w);
        $display("[%t ps][CPU ]: JAL rd[%d](%h), Jimm(%h)", $realtime, rd_id_w, (pc_r + 4), Jimm_w);
      end
      is_auipc_w: begin
        // $display("[%t ps][CPU ]: rd[%d] <- PC(%d) + Uimm(%h)", $realtime, rd_id_w, pc_r, Uimm_w);
        $display("[%t ps][CPU ]: AUIPC rd[%d], Uimm(%h)", $realtime, rd_id_w, Uimm_w);
      end
      is_lui_w: begin
        // $display("[%t ps][CPU ]: rd[%d] <- Uimm(%h)", $realtime, rd_id_w, Uimm_w);
        $display("[%t ps][CPU ]: LUI rd[%d], Uimm(%h)", $realtime, rd_id_w, Uimm_w);
      end
      is_load_w: begin
        // $display("[%t ps][CPU ]: rd[%d] <- MEM[rs1[%d] + Iimm(%h)]", $realtime, rd_id_w, rs1_id_w, Iimm_w);
        case (funct3_w)
          3'b000: $display("[%t ps][CPU ]: LB rd[%d], rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, Iimm_w);
          3'b001: $display("[%t ps][CPU ]: LH rd[%d], rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, Iimm_w);
          3'b010: $display("[%t ps][CPU ]: LW rd[%d], rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, Iimm_w);
          3'b100: $display("[%t ps][CPU ]: LBU rd[%d], rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, Iimm_w);
          3'b101: $display("[%t ps][CPU ]: LHU rd[%d], rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, Iimm_w);
          default: $display("[%t ps][CPU ]: Wrong Load, check funct3: rd[%d], rs1[%d](%h), Iimm(%h)", $realtime, rd_id_w, rs1_id_w, rs1_r, Iimm_w);
        endcase
      end
      is_store_w: begin
        // $display("[%t ps][CPU ]: MEM[rs1[%d] + Simm(%h)] <- rs2[%d]", $realtime, rs1_id_w, Simm_w, rs2_id_w);
        case (funct3_w)
          3'b000: $display("[%t ps][CPU ]: SB rs2[%d](%h), rs1[%d](%h), Simm(%h)", $realtime, rs2_id_w, rs2_r, rs1_id_w, rs1_r, Simm_w);
          3'b001: $display("[%t ps][CPU ]: SH rs2[%d](%h), rs1[%d](%h), Simm(%h)", $realtime, rs2_id_w, rs2_r, rs1_id_w, rs1_r, Simm_w);
          3'b010: $display("[%t ps][CPU ]: SW rs2[%d](%h), rs1[%d](%h), Simm(%h)", $realtime, rs2_id_w, rs2_r, rs1_id_w, rs1_r, Simm_w);
          default: $display("[%t ps][CPU ]: Wrong Store, check funct3: rs2[%d](%h), rs1[%d](%h), Iimm(%h)", $realtime, rs2_id_w, rs2_r, rs1_id_w, rs1_r, Simm_w);
        endcase
      end
      is_system_w: begin
        case (inst_r[20])
          1'b0: $display("[%t ps][CPU ]: ECALL(%h)", $realtime, inst_r);
          1'b1: begin
            $display("[%t ps][CPU ]: EBREAK(%h)", $realtime, inst_r);
            // $finish();
          end
          default: $display("[%t ps][CPU ]: System Instruction(%h)", $realtime, inst_r);
        endcase
      end
      default: $display("[%t ps][CPU ]: other instruction(%h)", $realtime, inst_r);
    endcase
  end
end

// ----------------------------------------------------------------------------
// ALU
// ----------------------------------------------------------------------------
// two types:
//     - Rtype: rd <- rs1 OP rs2 (is_alu_reg_w)
//     - Itype: rd <- rs1 OP Iimm (is_alu_imm_w)
wire [31:0] alu_in1_w = (
  (is_jal_w | is_jalr_w | is_auipc_w) ? pc_r : 
  (is_lui_w) ? 32'h0 : 
  rs1_r
);
wire [31:0] alu_in2_w = (
  (is_alu_reg_w | is_branch_w) ? rs2_r : 
  (is_auipc_w | is_lui_w) ? Uimm_w :
  (is_jal_w | is_jalr_w) ? 32'h4 :
  Iimm_w
);

wire [4:0] sh_amt_w = is_alu_reg_w ? rs2_r[4:0] : Iimm_w[4:0];

wire [31:0] alu_add_w = alu_in1_w + alu_in2_w;
wire [32:0] alu_sub_w = {1'b0, alu_in1_w} + {1'b1, ~alu_in2_w} + 33'b1;
wire [31:0] alu_ltu_w = {31'b0, alu_sub_w[32]};
wire [31:0] alu_lt_w = (alu_in1_w[31] ^ alu_in2_w[31]) ? {31'b0, alu_in1_w[31]} : alu_ltu_w;
wire [31:0] alu_xor_w = alu_in1_w ^ alu_in2_w;
wire [31:0] alu_or_w = alu_in1_w | alu_in2_w;
wire [31:0] alu_and_w = alu_in1_w & alu_in2_w;

// wire [31:0] signed_shift_right_w = $signed(alu_in1_w) >>> sh_amt_w; // SRA
// wire [31:0] unsigned_shift_right_w = alu_in1_w >> sh_amt_w;         // SRL
wire [32:0] alu_sra_w = $signed({(funct7_w[5] & alu_in1_w[31]), alu_in1_w}) >>> sh_amt_w;

reg [31:0] alu_out_w;
always @(*) begin
  case (funct3_w)
    // ADD or SUB
    // 3'b000: alu_out_w = (funct7_w[5] & inst_r[5]) ? (alu_in1_w - alu_in2_w) : (alu_in1_w + alu_in2_w);
    3'b000: alu_out_w = (funct7_w[5] & inst_r[5]) ? alu_sub_w[31:0] : alu_add_w;
    // left shift
    3'b001: alu_out_w = (alu_in1_w << sh_amt_w);
    // signed comparison (<)
    // 3'b010: alu_out_w = ($signed(alu_in1_w) < $signed(alu_in2_w));
    3'b010: alu_out_w = alu_lt_w;
    // unsigned comparison (<)
    // 3'b011: alu_out_w = (alu_in1_w < alu_in2_w);
    3'b011: alu_out_w = alu_ltu_w;
    // XOR
    3'b100: alu_out_w = alu_xor_w;
    // logical/arithmetic right shift
    3'b101: alu_out_w = alu_sra_w[31:0];
    // OR
    3'b110: alu_out_w = alu_or_w;
    // AND
    3'b111: alu_out_w = alu_and_w;
  endcase
end

reg [31:0] alu_out_r;
always @(posedge clk) begin
  if (rst) begin
    alu_out_r <= 32'b0;
  end
  else if (state_r == EXE) begin
    if (is_alu_reg_w | is_alu_imm_w) begin
      alu_out_r <= alu_out_w;
    end
    else begin
      alu_out_r <= alu_add_w;
    end
  end
  
end

// ----------------------------------------------------------------------------
// Branch
// ----------------------------------------------------------------------------
wire is_branch_ne_w = (|alu_xor_w);
wire is_branch_eq_w = (~is_branch_ne_w);
wire is_branch_lt_w = alu_lt_w;
wire is_branch_ge_w = (~alu_lt_w);
wire is_branch_ltu_w = alu_ltu_w;
wire is_branch_geu_w = (~alu_ltu_w);

reg is_branch_taken_w;
always @(*) begin
  case (funct3_w)
    // BEQ rs1, rs2, imm: if(rs1 == rs2) PC <- PC + Bimm
    // 3'b000: is_branch_taken_w = (rs1_r == rs2_r);
    3'b000: is_branch_taken_w = is_branch_eq_w;
    // BNE rs1, rs2, imm: if(rs1 != rs2) PC <- PC + Bimm
    // 3'b001: is_branch_taken_w = (rs1_r != rs2_r);
    3'b001: is_branch_taken_w = is_branch_ne_w;
    // BLT rs1, rs2, imm: if(rs1 < rs2) PC <- PC + Bimm (signed comparison)
    // 3'b100: is_branch_taken_w = ($signed(rs1_r) < $signed(rs2_r));
    3'b100: is_branch_taken_w = is_branch_lt_w;
    // BGE rs1, rs2, imm: if(rs1 >= rs2) PC <- PC + Bimm (signed comparison)
    // 3'b101: is_branch_taken_w = ($signed(rs1_r) >= $signed(rs2_r));
    3'b101: is_branch_taken_w = is_branch_ge_w;
    // BLTU rs1, rs2, imm: if(rs1 < rs2) PC <- PC + Bimm (unsigned comparison)
    // 3'b110: is_branch_taken_w = (rs1_r < rs2_r);
    3'b110: is_branch_taken_w = is_branch_ltu_w;
    // BGEU rs1, rs2, imm: if(rs1 >= rs2) PC <- PC + Bimm (unsigned comparison)
    // 3'b111: is_branch_taken_w = (rs1_r >= rs2_r);
    3'b111: is_branch_taken_w = is_branch_geu_w;
    // otherwise branch is not taken, `default` statement is necessary to avoid latch
    default: is_branch_taken_w = 1'b0;
  endcase
end

// wire [31:0] pc_plus_Bimm = pc_r + Bimm_w;

// ----------------------------------------------------------------------------
// Jump
// ----------------------------------------------------------------------------
// JAL rd, imm: rd <- PC + 4; PC <- PC + Jimm
// JALR rd, rs1, imm: rd <- PC + 4; PC <- rs1 + Iimm

// wire [31:0] pc_plus_4 = pc_r + 4;
// wire [31:0] pc_plus_4 = alu_out_w;
// wire [31:0] pc_plus_Jimm = pc_r + Jimm_w;
// wire [31:0] pc_plus_Uimm = pc_r + Uimm_w;
// wire [31:0] rs1_plus_Iimm = rs1_r + Iimm_w;

wire [31:0] next_pc_add1_w = is_jalr_w ? rs1_r : pc_r;
wire [31:0] next_pc_add2_w = (
  (is_branch_w & is_branch_taken_w) ? Bimm_w :
  (is_jal_w) ? Jimm_w :
  (is_jalr_w) ? Iimm_w :
  32'h4
);

// ----------------------------------------------------------------------------
// Generate Next PC
// ----------------------------------------------------------------------------
// wire [31:0] next_pc_w = (
//   (is_branch_w & is_branch_taken_w) ? pc_plus_Bimm :
//   (is_jal_w) ? pc_plus_Jimm :
//   (is_jalr_w) ? rs1_plus_Iimm :
//   pc_plus_4
// );
wire [31:0] next_pc_w = next_pc_add1_w + next_pc_add2_w;

reg [31:0] pc_r;
always @(posedge clk) begin
  if (rst) begin
    pc_r <= PC_BASE_ADDR;
  end
  else if (state_r == EXE) begin
    pc_r <= next_pc_w;
  end
end

// ----------------------------------------------------------------------------
// Load
// ----------------------------------------------------------------------------
wire [31:0] load_ori_addr_w = rs1_r + Iimm_w;
wire [31:0] load_word_addr_w = {load_ori_addr_w[31:2], 2'b0};

reg [31:0] load_ori_data_r;
always @(posedge clk) begin
  if (rst) begin
    load_ori_data_r <= 32'b0;
  end
  else if (state_r == MEM & is_load_w) begin
    load_ori_data_r <= mem_rdata_i;
  end
end

// convert mem_load_word to wb_load_word
wire is_load_store_byte_w = funct3_w[1:0] == 2'b00;
wire is_load_store_half_w = funct3_w[1:0] == 2'b01;
wire is_load_unsigned_w = funct3_w[2] == 1'b1;

wire [15:0] load_half_w = (
  load_ori_addr_w[1] ? load_ori_data_r[31:16] :
  load_ori_data_r[15:0]
);

wire [7:0] load_byte_w = (
  load_ori_addr_w[0] ? load_half_w[15:8] :
  load_half_w[7:0]
);

wire load_sign_w = (
  (~is_load_unsigned_w) & 
  (is_load_store_half_w ? load_half_w[15] : load_byte_w[7])
); 

wire [31:0] load_data_w = (
  is_load_store_half_w ? {{16{load_sign_w}}, load_half_w} :
  is_load_store_byte_w ? {{24{load_sign_w}}, load_byte_w} :
  load_ori_data_r
);

// ----------------------------------------------------------------------------
// Store
// ----------------------------------------------------------------------------
wire [31:0] store_ori_addr_w = rs1_r + Simm_w;
wire [31:0] store_word_addr_w = {store_ori_addr_w[31:2], 2'b0};

wire [31:0] store_byte_w = {4{rs2_r[7:0]}};
wire [31:0] store_half_w = {2{rs2_r[15:0]}};

wire [31:0] store_data_w = (
  is_load_store_byte_w ? store_byte_w :
  is_load_store_half_w ? store_half_w :
  rs2_r
);

wire [3:0] store_mask_w = (
  is_load_store_byte_w ? (
    store_ori_addr_w[0] ? (
      store_ori_addr_w[1] ? 4'b1000 : 4'b0010
    ) : (
      store_ori_addr_w[1] ? 4'b0100 : 4'b0001
    )
  ) :
  is_load_store_half_w ? (
    store_ori_addr_w[1] ? 4'b1100 : 4'b0011
  ) :
  4'b1111
);

// ----------------------------------------------------------------------------
// Write Back to rd
// ----------------------------------------------------------------------------
wire wb_en_w = (
  (state_r == WB) &
  (rd_id_w != 0) &
  (   
    is_alu_reg_w |
    is_alu_imm_w | 
    is_jal_w |
    is_jalr_w |
    is_auipc_w |
    is_lui_w |
    is_load_w
  )
);

wire [31:0] wb_data_w = is_load_w ? load_data_w : alu_out_r;

// ----------------------------------------------------------------------------
// Output Interface
// ----------------------------------------------------------------------------
assign mem_addr_o = (
  (state_r == EXE) ? (
    is_load_w ? load_word_addr_w :
    is_store_w ? store_word_addr_w :
    pc_r
  ) :
  pc_r
);

assign mem_rstrb_o = (
  (state_r == WB) |
  (state_r == EXE & is_load_w)
);

assign mem_wmask_o = (
  ((state_r == EXE) & (is_store_w)) ? store_mask_w :
  4'b0000
);

assign mem_wdata_o = store_data_w;

endmodule
